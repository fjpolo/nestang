// NES module to use rewind feature
// fjpolo, 01.2024

module NESrewind(
                    input i_clk,
                    input i_rst
                );

endmodule