`ifndef _wishbone_slaves_vh_
`define _wishbone_slaves_vh_

parameter WISHBONE_SLAVE_ADDRESS_TEST  = 1

`endif